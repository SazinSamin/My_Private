	module rtlfa32_4(s, cout, a, b, cin, clk);
		input [31:0] a,b;
		input cin, clk;
		output reg cout;
		output [31:0] s;
		reg [5:0] a1, a2, b1, b2, a22, b22, s1, s11, s111, s1111, s11111, s111111, s2, s22, s222, s2222, s22222, s1111111, s222222;
		reg [3:0] a3, a4, b3, b4, a33, a44, a333, a444, a4444, b333, b33, b44, b444, b4444;
		reg [3:0] s3, s33, s333, s3333, s4, s44, s4444, s33333, s444;
		reg c1, c2, c3, c4, c5, c6, ci;
		reg[3:0] a5,a55,a555,a5555,a55555,b5,b55,b555,b5555,b55555,s5,s55,s555;
		reg[3:0] a6,a66,a666,a6666,a66666,a666666,b6,b66,b666,b6666,b66666,b666666,s6,s66;
		reg[3:0] a7,a77,a777,a7777,a77777,a777777,a7777777,b7,b77,b777,b7777,b77777,b777777,b7777777,s7;


		always @ (posedge clk)
		        begin
		                a1<={a[5:0]};
		                a2<={a[11:6]};
		                a3<={a[15:12]};
		                a4<={a[19:16]};
		                a5<={a[23:20]};
				a6<={a[27:24]};
				a7<={a[31:28]};


		                b1<={b[5:0]};
		                b2<={b[11:6]};
		                b3<={b[15:12]};
		                b4<={b[19:16]};
		                b5<={b[23:20]};
				b6<={b[27:24]};
				b7<={b[31:28]};
		                ci<=cin;

		        end
		always @ (posedge clk)
		        begin
		          {c1,s1}<=a1+b1+ci;
		          a22<=a2;
			  b22<=b2;

		          a33<=a3;
		          a44<=a4;
		          b33<=b3;
		          b44<=b4;

		          a55<=a5;
		          b55<=b5;
			  a66<=a6;
		          b66<=b6;
			  
			  a77<=a7;
			  b77<=b7;


		        end
		always @ (posedge clk)
		        begin
		          s11<=s1;
		          {c2,s2}<=a22+b22+c1;
		          a333<=a33;
		          a444<=a44;
		          b333<=b33;
		          b444<=b44;

		          a555<=a55;
		          b555<=b55;

			  a666<=a66;
		          b666<=b66;
			  a777<=a77;
			  b777<=b77;


		        end

		always @ (posedge clk)
		        begin
		          s111<=s11;
		          s22<=s2;
			{c3,s3}<=a333+b333+c2;
		          a4444<=a444;
		          b4444<=b444;

		          a5555<=a555;
		          b5555<=b555;
			  a6666<=a666;
		          b6666<=b666;
			  a7777<=a777;
			  b7777<=b777;
		        end
		always @ (posedge clk)
		        begin
		          s1111<=s111;
		          s222<=s22;
		          s33<=s3;
		          {c4,s4}<=a4444+b4444+c3;

		          a55555<=a5555;
		          b55555<=b5555;
			  a66666<=a6666;
		          b66666<=b6666;
			  a77777<=a7777;
			  b77777<=b7777;


		        end

		     always @ (posedge clk)
		        begin
		          s11111<=s1111;
		          s2222<=s222;
		          s333<=s33;
		          s44<=s4;


		          {c5,s5}<=a55555+b55555+c4;
			
			  a666666<=a66666;
		          b666666<=b66666;
			  a777777<=a77777;
			  b777777<=b77777;



		        end


			 always @ (posedge clk)
					begin
					  s111111<=s11111;
					  s22222<=s2222;
		          		s3333<=s333;
		         		 s444<=s44;
					s55<=s5;
				{c6,s6}<=a666666+b666666+c5;
				
				a7777777<=a777777;
				b7777777<=b777777;
					  

					end
			
			always @ (posedge clk)
					begin
					  s1111111<=s111111;
					  s222222<=s22222;
		          		s33333<=s3333;
		         		 s4444<=s444;
					s555<=s55;
					s66<=s6;
				{cout,s7}<=a7777777+b7777777+c6;
					  
					end

			assign s={{s7[3:0]},{s66[3:0]},{s555[3:0]},{s4444[3:0]},{s33333[3:0]},{s222222[5:0]},{s1111111[5:0]}};

	endmodule
